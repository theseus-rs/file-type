<ColorDecisionList