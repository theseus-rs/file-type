<?xml version="1.0" encoding="ISO-8859-1"?>
<LENEX>
 <VERSION>