netcdf 